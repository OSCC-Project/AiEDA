//Generate the verilog at 2024-10-16T03:24:03
module gcd (
clk,
req_msg[31],
req_msg[30],
req_msg[29],
req_msg[28],
req_msg[27],
req_msg[26],
req_msg[25],
req_msg[24],
req_msg[23],
req_msg[22],
req_msg[21],
req_msg[20],
req_msg[19],
req_msg[18],
req_msg[17],
req_msg[16],
req_msg[15],
req_msg[14],
req_msg[13],
req_msg[12],
req_msg[11],
req_msg[10],
req_msg[9],
req_msg[8],
req_msg[7],
req_msg[6],
req_msg[5],
req_msg[4],
req_msg[3],
req_msg[2],
req_msg[1],
req_msg[0],
req_rdy,
req_val,
reset,
resp_msg[15],
resp_msg[14],
resp_msg[13],
resp_msg[12],
resp_msg[11],
resp_msg[10],
resp_msg[9],
resp_msg[8],
resp_msg[7],
resp_msg[6],
resp_msg[5],
resp_msg[4],
resp_msg[3],
resp_msg[2],
resp_msg[1],
resp_msg[0],
resp_rdy,
resp_val
);

input clk ;
input req_msg[31] ;
input req_msg[30] ;
input req_msg[29] ;
input req_msg[28] ;
input req_msg[27] ;
input req_msg[26] ;
input req_msg[25] ;
input req_msg[24] ;
input req_msg[23] ;
input req_msg[22] ;
input req_msg[21] ;
input req_msg[20] ;
input req_msg[19] ;
input req_msg[18] ;
input req_msg[17] ;
input req_msg[16] ;
input req_msg[15] ;
input req_msg[14] ;
input req_msg[13] ;
input req_msg[12] ;
input req_msg[11] ;
input req_msg[10] ;
input req_msg[9] ;
input req_msg[8] ;
input req_msg[7] ;
input req_msg[6] ;
input req_msg[5] ;
input req_msg[4] ;
input req_msg[3] ;
input req_msg[2] ;
input req_msg[1] ;
input req_msg[0] ;
output req_rdy ;
input req_val ;
input reset ;
output resp_msg[15] ;
output resp_msg[14] ;
output resp_msg[13] ;
output resp_msg[12] ;
output resp_msg[11] ;
output resp_msg[10] ;
output resp_msg[9] ;
output resp_msg[8] ;
output resp_msg[7] ;
output resp_msg[6] ;
output resp_msg[5] ;
output resp_msg[4] ;
output resp_msg[3] ;
output resp_msg[2] ;
output resp_msg[1] ;
output resp_msg[0] ;
input resp_rdy ;
output resp_val ;

wire clk ;
wire \req_msg[31] ;
wire \req_msg[30] ;
wire \req_msg[29] ;
wire \req_msg[28] ;
wire \req_msg[27] ;
wire \req_msg[26] ;
wire \req_msg[25] ;
wire \req_msg[24] ;
wire \req_msg[23] ;
wire \req_msg[22] ;
wire \req_msg[21] ;
wire \req_msg[20] ;
wire \req_msg[19] ;
wire \req_msg[18] ;
wire \req_msg[17] ;
wire \req_msg[16] ;
wire \req_msg[15] ;
wire \req_msg[14] ;
wire \req_msg[13] ;
wire \req_msg[12] ;
wire \req_msg[11] ;
wire \req_msg[10] ;
wire \req_msg[9] ;
wire \req_msg[8] ;
wire \req_msg[7] ;
wire \req_msg[6] ;
wire \req_msg[5] ;
wire \req_msg[4] ;
wire \req_msg[3] ;
wire \req_msg[2] ;
wire \req_msg[1] ;
wire \req_msg[0] ;
wire req_rdy ;
wire req_val ;
wire reset ;
wire \resp_msg[15] ;
wire \resp_msg[14] ;
wire \resp_msg[13] ;
wire \resp_msg[12] ;
wire \resp_msg[11] ;
wire \resp_msg[10] ;
wire \resp_msg[9] ;
wire \resp_msg[8] ;
wire \resp_msg[7] ;
wire \resp_msg[6] ;
wire \resp_msg[5] ;
wire \resp_msg[4] ;
wire \resp_msg[3] ;
wire \resp_msg[2] ;
wire \resp_msg[1] ;
wire \resp_msg[0] ;
wire resp_rdy ;
wire resp_val ;
wire ctrl_b_mux_sel_0_ ;
wire ctrl_b_reg_en_0_ ;
wire ctrl_a_reg_en_0_ ;
wire dpath_is_b_zero_0_ ;
wire dpath_is_a_lt_b_0_ ;
wire \ctrl_a_mux_sel[1] ;
wire \ctrl_a_mux_sel[0] ;
wire \ctrl/n1 ;
wire \ctrl/n2 ;
wire \ctrl/n3 ;
wire \ctrl/n4 ;
wire \ctrl/n5 ;
wire \ctrl/state_out[1] ;
wire \ctrl/state_out[0] ;
wire \ctrl/next_state__0[1] ;
wire \ctrl/next_state__0[0] ;
wire \ctrl/state/n1 ;
wire \dpath/n15 ;
wire \dpath/a_reg_out[15] ;
wire \dpath/a_reg_out[14] ;
wire \dpath/a_reg_out[13] ;
wire \dpath/a_reg_out[12] ;
wire \dpath/a_reg_out[11] ;
wire \dpath/a_reg_out[10] ;
wire \dpath/a_reg_out[9] ;
wire \dpath/a_reg_out[8] ;
wire \dpath/a_reg_out[7] ;
wire \dpath/a_reg_out[6] ;
wire \dpath/a_reg_out[5] ;
wire \dpath/a_reg_out[4] ;
wire \dpath/a_reg_out[3] ;
wire \dpath/a_reg_out[2] ;
wire \dpath/a_reg_out[1] ;
wire \dpath/a_reg_out[0] ;
wire \dpath/a_mux_out[15] ;
wire \dpath/a_mux_out[14] ;
wire \dpath/a_mux_out[13] ;
wire \dpath/a_mux_out[12] ;
wire \dpath/a_mux_out[11] ;
wire \dpath/a_mux_out[10] ;
wire \dpath/a_mux_out[9] ;
wire \dpath/a_mux_out[8] ;
wire \dpath/a_mux_out[7] ;
wire \dpath/a_mux_out[6] ;
wire \dpath/a_mux_out[5] ;
wire \dpath/a_mux_out[4] ;
wire \dpath/a_mux_out[3] ;
wire \dpath/a_mux_out[2] ;
wire \dpath/a_mux_out[1] ;
wire \dpath/a_mux_out[0] ;
wire \dpath/b_mux_out[15] ;
wire \dpath/b_mux_out[14] ;
wire \dpath/b_mux_out[13] ;
wire \dpath/b_mux_out[12] ;
wire \dpath/b_mux_out[11] ;
wire \dpath/b_mux_out[10] ;
wire \dpath/b_mux_out[9] ;
wire \dpath/b_mux_out[8] ;
wire \dpath/b_mux_out[7] ;
wire \dpath/b_mux_out[6] ;
wire \dpath/b_mux_out[5] ;
wire \dpath/b_mux_out[4] ;
wire \dpath/b_mux_out[3] ;
wire \dpath/b_mux_out[2] ;
wire \dpath/b_mux_out[1] ;
wire \dpath/b_mux_out[0] ;
wire \dpath/b_reg_out[15] ;
wire \dpath/b_reg_out[14] ;
wire \dpath/b_reg_out[13] ;
wire \dpath/b_reg_out[12] ;
wire \dpath/b_reg_out[11] ;
wire \dpath/b_reg_out[10] ;
wire \dpath/b_reg_out[9] ;
wire \dpath/b_reg_out[8] ;
wire \dpath/b_reg_out[7] ;
wire \dpath/b_reg_out[6] ;
wire \dpath/b_reg_out[5] ;
wire \dpath/b_reg_out[4] ;
wire \dpath/b_reg_out[3] ;
wire \dpath/b_reg_out[2] ;
wire \dpath/b_reg_out[1] ;
wire \dpath/b_reg_out[0] ;
wire \dpath/a_reg/n2 ;
wire \dpath/a_reg/n3 ;
wire \dpath/a_reg/n4 ;
wire \dpath/a_reg/n5 ;
wire \dpath/a_reg/n6 ;
wire \dpath/a_reg/n7 ;
wire \dpath/a_reg/n8 ;
wire \dpath/a_reg/n9 ;
wire \dpath/a_reg/n10 ;
wire \dpath/a_reg/n11 ;
wire \dpath/a_reg/n12 ;
wire \dpath/a_reg/n13 ;
wire \dpath/a_reg/n14 ;
wire \dpath/a_reg/n15 ;
wire \dpath/a_reg/n16 ;
wire \dpath/a_reg/n17 ;
wire \dpath/a_reg/n1 ;
wire \dpath/a_reg/n18 ;
wire \dpath/a_reg/n19 ;
wire \dpath/a_lt_b/n1 ;
wire \dpath/a_lt_b/n2 ;
wire \dpath/a_lt_b/n3 ;
wire \dpath/a_lt_b/n4 ;
wire \dpath/a_lt_b/n5 ;
wire \dpath/a_lt_b/n6 ;
wire \dpath/a_lt_b/n7 ;
wire \dpath/a_lt_b/n8 ;
wire \dpath/a_lt_b/n9 ;
wire \dpath/a_lt_b/n10 ;
wire \dpath/a_lt_b/n11 ;
wire \dpath/a_lt_b/n12 ;
wire \dpath/a_lt_b/n13 ;
wire \dpath/a_lt_b/n14 ;
wire \dpath/a_lt_b/n15 ;
wire \dpath/a_lt_b/n16 ;
wire \dpath/a_lt_b/n17 ;
wire \dpath/a_lt_b/n18 ;
wire \dpath/a_lt_b/n19 ;
wire \dpath/a_lt_b/n20 ;
wire \dpath/a_lt_b/n21 ;
wire \dpath/a_lt_b/n22 ;
wire \dpath/a_lt_b/n23 ;
wire \dpath/a_lt_b/n24 ;
wire \dpath/a_lt_b/n25 ;
wire \dpath/a_lt_b/n26 ;
wire \dpath/a_lt_b/n27 ;
wire \dpath/a_lt_b/n28 ;
wire \dpath/a_lt_b/n29 ;
wire \dpath/a_lt_b/n30 ;
wire \dpath/a_lt_b/n31 ;
wire \dpath/a_lt_b/n32 ;
wire \dpath/a_lt_b/n33 ;
wire \dpath/a_lt_b/n34 ;
wire \dpath/a_lt_b/n35 ;
wire \dpath/a_lt_b/n36 ;
wire \dpath/a_lt_b/n37 ;
wire \dpath/b_zero/n1 ;
wire \dpath/b_zero/n2 ;
wire \dpath/b_zero/n3 ;
wire \dpath/b_zero/n4 ;
wire \dpath/a_mux/n1 ;
wire \dpath/a_mux/n2 ;
wire \dpath/a_mux/n3 ;
wire \dpath/a_mux/n4 ;
wire \dpath/a_mux/n5 ;
wire \dpath/a_mux/n6 ;
wire \dpath/a_mux/n7 ;
wire \dpath/a_mux/n8 ;
wire \dpath/a_mux/n9 ;
wire \dpath/a_mux/n10 ;
wire \dpath/a_mux/n11 ;
wire \dpath/a_mux/n12 ;
wire \dpath/a_mux/n13 ;
wire \dpath/a_mux/n14 ;
wire \dpath/a_mux/n15 ;
wire \dpath/a_mux/n16 ;
wire \dpath/a_mux/n17 ;
wire \dpath/a_mux/n18 ;
wire \dpath/b_mux/n1 ;
wire \dpath/sub/n45 ;
wire \dpath/sub/n46 ;
wire \dpath/sub/n47 ;
wire \dpath/sub/n48 ;
wire \dpath/sub/n49 ;
wire \dpath/sub/n50 ;
wire \dpath/sub/n1 ;
wire \dpath/sub/n3 ;
wire \dpath/sub/n5 ;
wire \dpath/sub/n7 ;
wire \dpath/sub/n9 ;
wire \dpath/sub/n11 ;
wire \dpath/sub/n13 ;
wire \dpath/sub/n14 ;
wire \dpath/sub/n15 ;
wire \dpath/sub/n16 ;
wire \dpath/sub/n17 ;
wire \dpath/sub/n18 ;
wire \dpath/sub/n19 ;
wire \dpath/sub/n20 ;
wire \dpath/sub/n21 ;
wire \dpath/sub/n22 ;
wire \dpath/sub/n23 ;
wire \dpath/sub/n24 ;
wire \dpath/sub/n25 ;
wire \dpath/sub/n26 ;
wire \dpath/sub/n27 ;
wire \dpath/sub/n28 ;
wire \dpath/sub/n29 ;
wire \dpath/sub/n30 ;
wire \dpath/sub/n31 ;
wire \dpath/sub/n32 ;
wire \dpath/sub/n33 ;
wire \dpath/sub/n34 ;
wire \dpath/sub/n35 ;
wire \dpath/sub/n36 ;
wire \dpath/sub/n37 ;
wire \dpath/sub/n38 ;
wire \dpath/sub/n39 ;
wire \dpath/sub/n40 ;
wire \dpath/sub/n41 ;
wire \dpath/sub/n42 ;
wire \dpath/sub/n43 ;
wire \dpath/sub/n44 ;
wire \dpath/b_reg/n2 ;
wire \dpath/b_reg/n3 ;
wire \dpath/b_reg/n4 ;
wire \dpath/b_reg/n5 ;
wire \dpath/b_reg/n6 ;
wire \dpath/b_reg/n7 ;
wire \dpath/b_reg/n8 ;
wire \dpath/b_reg/n9 ;
wire \dpath/b_reg/n10 ;
wire \dpath/b_reg/n11 ;
wire \dpath/b_reg/n12 ;
wire \dpath/b_reg/n13 ;
wire \dpath/b_reg/n14 ;
wire \dpath/b_reg/n15 ;
wire \dpath/b_reg/n16 ;
wire \dpath/b_reg/n17 ;
wire \dpath/b_reg/n1 ;
wire clk_0 ;
wire clk_1 ;

assign \req_msg[31] = req_msg[31] ;
assign \req_msg[30] = req_msg[30] ;
assign \req_msg[29] = req_msg[29] ;
assign \req_msg[28] = req_msg[28] ;
assign \req_msg[27] = req_msg[27] ;
assign \req_msg[26] = req_msg[26] ;
assign \req_msg[25] = req_msg[25] ;
assign \req_msg[24] = req_msg[24] ;
assign \req_msg[23] = req_msg[23] ;
assign \req_msg[22] = req_msg[22] ;
assign \req_msg[21] = req_msg[21] ;
assign \req_msg[20] = req_msg[20] ;
assign \req_msg[19] = req_msg[19] ;
assign \req_msg[18] = req_msg[18] ;
assign \req_msg[17] = req_msg[17] ;
assign \req_msg[16] = req_msg[16] ;
assign \req_msg[15] = req_msg[15] ;
assign \req_msg[14] = req_msg[14] ;
assign \req_msg[13] = req_msg[13] ;
assign \req_msg[12] = req_msg[12] ;
assign \req_msg[11] = req_msg[11] ;
assign \req_msg[10] = req_msg[10] ;
assign \req_msg[9] = req_msg[9] ;
assign \req_msg[8] = req_msg[8] ;
assign \req_msg[7] = req_msg[7] ;
assign \req_msg[6] = req_msg[6] ;
assign \req_msg[5] = req_msg[5] ;
assign \req_msg[4] = req_msg[4] ;
assign \req_msg[3] = req_msg[3] ;
assign \req_msg[2] = req_msg[2] ;
assign \req_msg[1] = req_msg[1] ;
assign \req_msg[0] = req_msg[0] ;
assign resp_msg[15] = \resp_msg[15] ;
assign resp_msg[14] = \resp_msg[14] ;
assign resp_msg[13] = \resp_msg[13] ;
assign resp_msg[12] = \resp_msg[12] ;
assign resp_msg[11] = \resp_msg[11] ;
assign resp_msg[10] = \resp_msg[10] ;
assign resp_msg[9] = \resp_msg[9] ;
assign resp_msg[8] = \resp_msg[8] ;
assign resp_msg[7] = \resp_msg[7] ;
assign resp_msg[6] = \resp_msg[6] ;
assign resp_msg[5] = \resp_msg[5] ;
assign resp_msg[4] = \resp_msg[4] ;
assign resp_msg[3] = \resp_msg[3] ;
assign resp_msg[2] = \resp_msg[2] ;
assign resp_msg[1] = \resp_msg[1] ;
assign resp_msg[0] = \resp_msg[0] ;

AOI21D1BWP40P140 \ctrl/U3 ( .ZN(ctrl_b_reg_en_0_ ), .B(\ctrl/state_out[1] ), .A2(\ctrl/n3 ), .A1(\ctrl/state_out[0] ) );
INVD1BWP40P140 \ctrl/U4 ( .ZN(ctrl_a_reg_en_0_ ), .I(\ctrl/state_out[1] ) );
NR2D1BWP40P140 \ctrl/U5 ( .ZN(ctrl_b_mux_sel_0_ ), .A2(\ctrl/state_out[0] ), .A1(\ctrl/state_out[1] ) );
BUFFD3BWP40P140 \ctrl/U7 ( .Z(req_rdy ), .I(ctrl_b_mux_sel_0_ ) );
ND2D1BWP40P140 \ctrl/U8 ( .ZN(\ctrl/n2 ), .A2(\ctrl/state_out[0] ), .A1(ctrl_a_reg_en_0_ ) );
NR2D1BWP40P140 \ctrl/U9 ( .ZN(\ctrl_a_mux_sel[0] ), .A2(\ctrl/n2 ), .A1(dpath_is_a_lt_b_0_ ) );
AOI21D1BWP40P140 \ctrl/U10 ( .ZN(\ctrl/n1 ), .B(\ctrl/state_out[0] ), .A2(ctrl_a_reg_en_0_ ), .A1(req_val ) );
AOI21D1BWP40P140 \ctrl/U11 ( .ZN(\ctrl/next_state__0[0] ), .B(\ctrl/n1 ), .A2(\ctrl_a_mux_sel[0] ), .A1(dpath_is_b_zero_0_ ) );
INVD1BWP40P140 \ctrl/U12 ( .ZN(\ctrl/n3 ), .I(dpath_is_a_lt_b_0_ ) );
NR2D1BWP40P140 \ctrl/U13 ( .ZN(\ctrl_a_mux_sel[1] ), .A2(\ctrl/n2 ), .A1(\ctrl/n3 ) );
INVD1BWP40P140 \ctrl/U14 ( .ZN(\ctrl/n5 ), .I(\ctrl/state_out[0] ) );
ND2D1BWP40P140 \ctrl/U15 ( .ZN(\ctrl/n4 ), .A2(dpath_is_b_zero_0_ ), .A1(\ctrl_a_mux_sel[0] ) );
AOI22D1BWP40P140 \ctrl/U16 ( .ZN(\ctrl/next_state__0[1] ), .B2(ctrl_a_reg_en_0_ ), .B1(\ctrl/n4 ), .A2(resp_rdy ), .A1(\ctrl/n5 ) );
DFKCNQD1BWP40P140 \ctrl/state/out_reg_1_ ( .Q(\ctrl/state_out[1] ), .D(\ctrl/next_state__0[1] ), .CP(clk_0 ), .CN(\ctrl/state/n1 ) );
DFKCNQD1BWP40P140 \ctrl/state/out_reg_0_ ( .Q(\ctrl/state_out[0] ), .D(\ctrl/next_state__0[0] ), .CP(clk_0 ), .CN(\ctrl/state/n1 ) );
INVD1BWP40P140 \ctrl/state/U3 ( .ZN(\ctrl/state/n1 ), .I(reset ) );
NR2OPTPAD4BWP40P140 \ctrl/U6 ( .ZN(resp_val ), .A2(ctrl_a_reg_en_0_ ), .A1(\ctrl/state_out[0] ) );
BUFFD3BWP40P140 \dpath/U1 ( .Z(\resp_msg[0] ), .I(\dpath/n15 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_15_ ( .Q(\dpath/a_reg_out[15] ), .D(\dpath/a_reg/n17 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_14_ ( .Q(\dpath/a_reg_out[14] ), .D(\dpath/a_reg/n16 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_13_ ( .Q(\dpath/a_reg_out[13] ), .D(\dpath/a_reg/n15 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_12_ ( .Q(\dpath/a_reg_out[12] ), .D(\dpath/a_reg/n14 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_11_ ( .Q(\dpath/a_reg_out[11] ), .D(\dpath/a_reg/n13 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_9_ ( .Q(\dpath/a_reg_out[9] ), .D(\dpath/a_reg/n11 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_8_ ( .Q(\dpath/a_reg_out[8] ), .D(\dpath/a_reg/n10 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_7_ ( .Q(\dpath/a_reg_out[7] ), .D(\dpath/a_reg/n9 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_6_ ( .Q(\dpath/a_reg_out[6] ), .D(\dpath/a_reg/n8 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_5_ ( .Q(\dpath/a_reg_out[5] ), .D(\dpath/a_reg/n7 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_4_ ( .Q(\dpath/a_reg_out[4] ), .D(\dpath/a_reg/n6 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_3_ ( .Q(\dpath/a_reg_out[3] ), .D(\dpath/a_reg/n5 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_2_ ( .Q(\dpath/a_reg_out[2] ), .D(\dpath/a_reg/n4 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_0_ ( .Q(\dpath/a_reg_out[0] ), .D(\dpath/a_reg/n2 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/a_reg/out_reg_1_ ( .Q(\dpath/a_reg_out[1] ), .D(\dpath/a_reg/n3 ), .CP(clk_0 ) );
MOAI22D1BWP40P140 \dpath/a_reg/U2 ( .ZN(\dpath/a_reg/n16 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[14] ), .A2(\dpath/a_reg/n1 ), .A1(\dpath/a_reg/n18 ) );
INVD1BWP40P140 \dpath/a_reg/U3 ( .ZN(\dpath/a_reg/n1 ), .I(\dpath/a_mux_out[14] ) );
INVD1BWP40P140 \dpath/a_reg/U4 ( .ZN(\dpath/a_reg/n18 ), .I(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U5 ( .Z(\dpath/a_reg/n17 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[15] ), .A2(\dpath/a_mux_out[15] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U6 ( .Z(\dpath/a_reg/n15 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[13] ), .A2(\dpath/a_mux_out[13] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U7 ( .Z(\dpath/a_reg/n14 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[12] ), .A2(\dpath/a_mux_out[12] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U8 ( .Z(\dpath/a_reg/n13 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[11] ), .A2(\dpath/a_mux_out[11] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U9 ( .Z(\dpath/a_reg/n12 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[10] ), .A2(\dpath/a_mux_out[10] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U10 ( .Z(\dpath/a_reg/n11 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[9] ), .A2(\dpath/a_mux_out[9] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U11 ( .Z(\dpath/a_reg/n10 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[8] ), .A2(\dpath/a_mux_out[8] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U12 ( .Z(\dpath/a_reg/n9 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[7] ), .A2(\dpath/a_mux_out[7] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U13 ( .Z(\dpath/a_reg/n8 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[6] ), .A2(\dpath/a_mux_out[6] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U14 ( .Z(\dpath/a_reg/n7 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[5] ), .A2(\dpath/a_mux_out[5] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U15 ( .Z(\dpath/a_reg/n6 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[4] ), .A2(\dpath/a_mux_out[4] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U16 ( .Z(\dpath/a_reg/n5 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[3] ), .A2(\dpath/a_mux_out[3] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U17 ( .Z(\dpath/a_reg/n4 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[2] ), .A2(\dpath/a_mux_out[2] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U18 ( .Z(\dpath/a_reg/n3 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[1] ), .A2(\dpath/a_mux_out[1] ), .A1(ctrl_a_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/a_reg/U19 ( .Z(\dpath/a_reg/n2 ), .B2(\dpath/a_reg/n18 ), .B1(\dpath/a_reg_out[0] ), .A2(\dpath/a_mux_out[0] ), .A1(ctrl_a_reg_en_0_ ) );
DFKCNQD1BWP40P140 \dpath/a_reg/out_reg_10_ ( .Q(\dpath/a_reg_out[10] ), .D(\dpath/a_reg/n19 ), .CP(clk_1 ), .CN(\dpath/a_reg/n12 ) );
TIEHBWP40P140LVT \dpath/a_reg/U20 ( .Z(\dpath/a_reg/n19 ) );
INVD1BWP40P140 \dpath/a_lt_b/U1 ( .ZN(\dpath/a_lt_b/n37 ), .I(\dpath/a_reg_out[15] ) );
INVD1BWP40P140 \dpath/a_lt_b/U2 ( .ZN(\dpath/a_lt_b/n32 ), .I(\dpath/a_reg_out[13] ) );
INVD1BWP40P140 \dpath/a_lt_b/U3 ( .ZN(\dpath/a_lt_b/n27 ), .I(\dpath/a_reg_out[11] ) );
INVD1BWP40P140 \dpath/a_lt_b/U4 ( .ZN(\dpath/a_lt_b/n24 ), .I(\dpath/a_reg_out[10] ) );
INVD1BWP40P140 \dpath/a_lt_b/U5 ( .ZN(\dpath/a_lt_b/n18 ), .I(\dpath/b_reg_out[9] ) );
MAOI22D1BWP40P140 \dpath/a_lt_b/U6 ( .ZN(\dpath/a_lt_b/n23 ), .B2(\dpath/b_reg_out[10] ), .B1(\dpath/a_lt_b/n24 ), .A2(\dpath/a_lt_b/n18 ), .A1(\dpath/a_reg_out[9] ) );
INVD1BWP40P140 \dpath/a_lt_b/U7 ( .ZN(\dpath/a_lt_b/n10 ), .I(\dpath/a_reg_out[5] ) );
INVD1BWP40P140 \dpath/a_lt_b/U8 ( .ZN(\dpath/a_lt_b/n4 ), .I(\dpath/b_reg_out[3] ) );
INVD1BWP40P140 \dpath/a_lt_b/U9 ( .ZN(\dpath/a_lt_b/n12 ), .I(\dpath/b_reg_out[4] ) );
AOI22D1BWP40P140 \dpath/a_lt_b/U10 ( .ZN(\dpath/a_lt_b/n9 ), .B2(\dpath/a_lt_b/n12 ), .B1(\dpath/a_reg_out[4] ), .A2(\dpath/a_lt_b/n4 ), .A1(\dpath/a_reg_out[3] ) );
INVD1BWP40P140 \dpath/a_lt_b/U11 ( .ZN(\dpath/a_lt_b/n3 ), .I(\dpath/b_reg_out[1] ) );
INVD1BWP40P140 \dpath/a_lt_b/U12 ( .ZN(\dpath/a_lt_b/n1 ), .I(\dpath/b_reg_out[0] ) );
OAI22D1BWP40P140 \dpath/a_lt_b/U13 ( .ZN(\dpath/a_lt_b/n2 ), .B2(\dpath/a_reg_out[0] ), .B1(\dpath/a_lt_b/n1 ), .A2(\dpath/a_lt_b/n3 ), .A1(\dpath/a_reg_out[1] ) );
IOA21D1BWP40P140 \dpath/a_lt_b/U14 ( .ZN(\dpath/a_lt_b/n7 ), .B(\dpath/a_lt_b/n2 ), .A2(\dpath/a_reg_out[1] ), .A1(\dpath/a_lt_b/n3 ) );
OR2D1BWP40P140 \dpath/a_lt_b/U15 ( .Z(\dpath/a_lt_b/n6 ), .A2(\dpath/a_lt_b/n4 ), .A1(\dpath/a_reg_out[3] ) );
IOA21D1BWP40P140 \dpath/a_lt_b/U16 ( .ZN(\dpath/a_lt_b/n5 ), .B(\dpath/b_reg_out[2] ), .A2(\dpath/a_reg_out[2] ), .A1(\dpath/a_lt_b/n7 ) );
OAI211D1BWP40P140 \dpath/a_lt_b/U17 ( .ZN(\dpath/a_lt_b/n8 ), .C(\dpath/a_lt_b/n5 ), .B(\dpath/a_lt_b/n6 ), .A2(\dpath/a_reg_out[2] ), .A1(\dpath/a_lt_b/n7 ) );
AOI22D1BWP40P140 \dpath/a_lt_b/U18 ( .ZN(\dpath/a_lt_b/n13 ), .B2(\dpath/a_lt_b/n8 ), .B1(\dpath/a_lt_b/n9 ), .A2(\dpath/a_lt_b/n10 ), .A1(\dpath/b_reg_out[5] ) );
INVD1BWP40P140 \dpath/a_lt_b/U19 ( .ZN(\dpath/a_lt_b/n14 ), .I(\dpath/b_reg_out[6] ) );
MOAI22D1BWP40P140 \dpath/a_lt_b/U20 ( .ZN(\dpath/a_lt_b/n11 ), .B2(\dpath/a_reg_out[6] ), .B1(\dpath/a_lt_b/n14 ), .A2(\dpath/a_lt_b/n10 ), .A1(\dpath/b_reg_out[5] ) );
AOI221D1BWP40P140 \dpath/a_lt_b/U21 ( .ZN(\dpath/a_lt_b/n17 ), .C(\dpath/a_lt_b/n11 ), .B2(\dpath/a_lt_b/n13 ), .B1(\dpath/a_lt_b/n12 ), .A2(\dpath/a_lt_b/n13 ), .A1(\dpath/a_reg_out[4] ) );
INVD1BWP40P140 \dpath/a_lt_b/U22 ( .ZN(\dpath/a_lt_b/n15 ), .I(\dpath/a_reg_out[7] ) );
MOAI22D1BWP40P140 \dpath/a_lt_b/U23 ( .ZN(\dpath/a_lt_b/n16 ), .B2(\dpath/b_reg_out[7] ), .B1(\dpath/a_lt_b/n15 ), .A2(\dpath/a_lt_b/n14 ), .A1(\dpath/a_reg_out[6] ) );
OAI22D1BWP40P140 \dpath/a_lt_b/U24 ( .ZN(\dpath/a_lt_b/n21 ), .B2(\dpath/a_lt_b/n15 ), .B1(\dpath/b_reg_out[7] ), .A2(\dpath/a_lt_b/n16 ), .A1(\dpath/a_lt_b/n17 ) );
OR2D1BWP40P140 \dpath/a_lt_b/U25 ( .Z(\dpath/a_lt_b/n20 ), .A2(\dpath/a_lt_b/n18 ), .A1(\dpath/a_reg_out[9] ) );
IOA21D1BWP40P140 \dpath/a_lt_b/U26 ( .ZN(\dpath/a_lt_b/n19 ), .B(\dpath/b_reg_out[8] ), .A2(\dpath/a_reg_out[8] ), .A1(\dpath/a_lt_b/n21 ) );
OAI211D1BWP40P140 \dpath/a_lt_b/U27 ( .ZN(\dpath/a_lt_b/n22 ), .C(\dpath/a_lt_b/n19 ), .B(\dpath/a_lt_b/n20 ), .A2(\dpath/a_reg_out[8] ), .A1(\dpath/a_lt_b/n21 ) );
AOI22D1BWP40P140 \dpath/a_lt_b/U28 ( .ZN(\dpath/a_lt_b/n25 ), .B2(\dpath/a_lt_b/n22 ), .B1(\dpath/a_lt_b/n23 ), .A2(\dpath/a_lt_b/n24 ), .A1(\dpath/b_reg_out[10] ) );
IOA21D1BWP40P140 \dpath/a_lt_b/U29 ( .ZN(\dpath/a_lt_b/n26 ), .B(\dpath/a_lt_b/n25 ), .A2(\dpath/b_reg_out[11] ), .A1(\dpath/a_lt_b/n27 ) );
OAI21D1BWP40P140 \dpath/a_lt_b/U30 ( .ZN(\dpath/a_lt_b/n30 ), .B(\dpath/a_lt_b/n26 ), .A2(\dpath/a_lt_b/n27 ), .A1(\dpath/b_reg_out[11] ) );
ND2D1BWP40P140 \dpath/a_lt_b/U31 ( .ZN(\dpath/a_lt_b/n29 ), .A2(\dpath/b_reg_out[13] ), .A1(\dpath/a_lt_b/n32 ) );
IOA21D1BWP40P140 \dpath/a_lt_b/U32 ( .ZN(\dpath/a_lt_b/n28 ), .B(\dpath/b_reg_out[12] ), .A2(\dpath/a_reg_out[12] ), .A1(\dpath/a_lt_b/n30 ) );
OAI211D1BWP40P140 \dpath/a_lt_b/U33 ( .ZN(\dpath/a_lt_b/n31 ), .C(\dpath/a_lt_b/n28 ), .B(\dpath/a_lt_b/n29 ), .A2(\dpath/a_reg_out[12] ), .A1(\dpath/a_lt_b/n30 ) );
OAI21D1BWP40P140 \dpath/a_lt_b/U34 ( .ZN(\dpath/a_lt_b/n35 ), .B(\dpath/a_lt_b/n31 ), .A2(\dpath/a_lt_b/n32 ), .A1(\dpath/b_reg_out[13] ) );
ND2D1BWP40P140 \dpath/a_lt_b/U35 ( .ZN(\dpath/a_lt_b/n34 ), .A2(\dpath/b_reg_out[15] ), .A1(\dpath/a_lt_b/n37 ) );
IOA21D1BWP40P140 \dpath/a_lt_b/U36 ( .ZN(\dpath/a_lt_b/n33 ), .B(\dpath/b_reg_out[14] ), .A2(\dpath/a_reg_out[14] ), .A1(\dpath/a_lt_b/n35 ) );
OAI211D1BWP40P140 \dpath/a_lt_b/U37 ( .ZN(\dpath/a_lt_b/n36 ), .C(\dpath/a_lt_b/n33 ), .B(\dpath/a_lt_b/n34 ), .A2(\dpath/a_reg_out[14] ), .A1(\dpath/a_lt_b/n35 ) );
OA21D1BWP40P140 \dpath/a_lt_b/U38 ( .Z(dpath_is_a_lt_b_0_ ), .B(\dpath/a_lt_b/n36 ), .A2(\dpath/a_lt_b/n37 ), .A1(\dpath/b_reg_out[15] ) );
OR4D1BWP40P140 \dpath/b_zero/U1 ( .Z(\dpath/b_zero/n4 ), .A4(\dpath/b_reg_out[15] ), .A3(\dpath/b_reg_out[14] ), .A2(\dpath/b_reg_out[13] ), .A1(\dpath/b_reg_out[12] ) );
OR4D1BWP40P140 \dpath/b_zero/U2 ( .Z(\dpath/b_zero/n3 ), .A4(\dpath/b_reg_out[11] ), .A3(\dpath/b_reg_out[10] ), .A2(\dpath/b_reg_out[9] ), .A1(\dpath/b_reg_out[8] ) );
OR4D1BWP40P140 \dpath/b_zero/U3 ( .Z(\dpath/b_zero/n2 ), .A4(\dpath/b_reg_out[7] ), .A3(\dpath/b_reg_out[6] ), .A2(\dpath/b_reg_out[5] ), .A1(\dpath/b_reg_out[4] ) );
OR4D1BWP40P140 \dpath/b_zero/U4 ( .Z(\dpath/b_zero/n1 ), .A4(\dpath/b_reg_out[3] ), .A3(\dpath/b_reg_out[2] ), .A2(\dpath/b_reg_out[1] ), .A1(\dpath/b_reg_out[0] ) );
NR4D1BWP40P140 \dpath/b_zero/U5 ( .ZN(dpath_is_b_zero_0_ ), .A4(\dpath/b_zero/n1 ), .A3(\dpath/b_zero/n2 ), .A2(\dpath/b_zero/n3 ), .A1(\dpath/b_zero/n4 ) );
IOA21D1BWP40P140 \dpath/a_mux/U1 ( .ZN(\dpath/a_mux_out[14] ), .B(\dpath/a_mux/n1 ), .A2(\resp_msg[14] ), .A1(\dpath/a_mux/n18 ) );
INR2D1BWP40P140 \dpath/a_mux/U2 ( .ZN(\dpath/a_mux/n18 ), .B1(\ctrl_a_mux_sel[1] ), .A1(\ctrl_a_mux_sel[0] ) );
NR2D1BWP40P140 \dpath/a_mux/U3 ( .ZN(\dpath/a_mux/n16 ), .A2(\ctrl_a_mux_sel[0] ), .A1(\ctrl_a_mux_sel[1] ) );
AOI22D1BWP40P140 \dpath/a_mux/U4 ( .ZN(\dpath/a_mux/n1 ), .B2(\req_msg[30] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[14] ), .A1(\ctrl_a_mux_sel[1] ) );
AOI22D1BWP40P140 \dpath/a_mux/U5 ( .ZN(\dpath/a_mux/n2 ), .B2(\req_msg[27] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[11] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U6 ( .ZN(\dpath/a_mux_out[11] ), .B(\dpath/a_mux/n2 ), .A2(\resp_msg[11] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U7 ( .ZN(\dpath/a_mux/n3 ), .B2(\req_msg[17] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[1] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U8 ( .ZN(\dpath/a_mux_out[1] ), .B(\dpath/a_mux/n3 ), .A2(\resp_msg[1] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U9 ( .ZN(\dpath/a_mux/n4 ), .B2(\req_msg[24] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[8] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U10 ( .ZN(\dpath/a_mux_out[8] ), .B(\dpath/a_mux/n4 ), .A2(\resp_msg[8] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U11 ( .ZN(\dpath/a_mux/n5 ), .B2(\req_msg[16] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[0] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U12 ( .ZN(\dpath/a_mux_out[0] ), .B(\dpath/a_mux/n5 ), .A2(\resp_msg[0] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U13 ( .ZN(\dpath/a_mux/n6 ), .B2(\req_msg[19] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[3] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U14 ( .ZN(\dpath/a_mux_out[3] ), .B(\dpath/a_mux/n6 ), .A2(\resp_msg[3] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U15 ( .ZN(\dpath/a_mux/n7 ), .B2(\req_msg[20] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[4] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U16 ( .ZN(\dpath/a_mux_out[4] ), .B(\dpath/a_mux/n7 ), .A2(\resp_msg[4] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U17 ( .ZN(\dpath/a_mux/n8 ), .B2(\req_msg[18] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[2] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U18 ( .ZN(\dpath/a_mux_out[2] ), .B(\dpath/a_mux/n8 ), .A2(\resp_msg[2] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U19 ( .ZN(\dpath/a_mux/n9 ), .B2(\req_msg[23] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[7] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U20 ( .ZN(\dpath/a_mux_out[7] ), .B(\dpath/a_mux/n9 ), .A2(\resp_msg[7] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U21 ( .ZN(\dpath/a_mux/n10 ), .B2(\req_msg[28] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[12] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U22 ( .ZN(\dpath/a_mux_out[12] ), .B(\dpath/a_mux/n10 ), .A2(\resp_msg[12] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U23 ( .ZN(\dpath/a_mux/n11 ), .B2(\req_msg[29] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[13] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U24 ( .ZN(\dpath/a_mux_out[13] ), .B(\dpath/a_mux/n11 ), .A2(\resp_msg[13] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U25 ( .ZN(\dpath/a_mux/n12 ), .B2(\req_msg[31] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[15] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U26 ( .ZN(\dpath/a_mux_out[15] ), .B(\dpath/a_mux/n12 ), .A2(\resp_msg[15] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U27 ( .ZN(\dpath/a_mux/n13 ), .B2(\req_msg[21] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[5] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U28 ( .ZN(\dpath/a_mux_out[5] ), .B(\dpath/a_mux/n13 ), .A2(\resp_msg[5] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U29 ( .ZN(\dpath/a_mux/n14 ), .B2(\req_msg[22] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[6] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U30 ( .ZN(\dpath/a_mux_out[6] ), .B(\dpath/a_mux/n14 ), .A2(\resp_msg[6] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U31 ( .ZN(\dpath/a_mux/n15 ), .B2(\req_msg[25] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[9] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U32 ( .ZN(\dpath/a_mux_out[9] ), .B(\dpath/a_mux/n15 ), .A2(\resp_msg[9] ), .A1(\dpath/a_mux/n18 ) );
AOI22D1BWP40P140 \dpath/a_mux/U33 ( .ZN(\dpath/a_mux/n17 ), .B2(\req_msg[26] ), .B1(\dpath/a_mux/n16 ), .A2(\dpath/b_reg_out[10] ), .A1(\ctrl_a_mux_sel[1] ) );
IOA21D1BWP40P140 \dpath/a_mux/U34 ( .ZN(\dpath/a_mux_out[10] ), .B(\dpath/a_mux/n17 ), .A2(\resp_msg[10] ), .A1(\dpath/a_mux/n18 ) );
INVD1BWP40P140 \dpath/b_mux/U1 ( .ZN(\dpath/b_mux/n1 ), .I(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U2 ( .Z(\dpath/b_mux_out[0] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[0] ), .A2(\req_msg[0] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U3 ( .Z(\dpath/b_mux_out[1] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[1] ), .A2(\req_msg[1] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U4 ( .Z(\dpath/b_mux_out[2] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[2] ), .A2(\req_msg[2] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U5 ( .Z(\dpath/b_mux_out[3] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[3] ), .A2(\req_msg[3] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U6 ( .Z(\dpath/b_mux_out[4] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[4] ), .A2(\req_msg[4] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U7 ( .Z(\dpath/b_mux_out[5] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[5] ), .A2(\req_msg[5] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U8 ( .Z(\dpath/b_mux_out[6] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[6] ), .A2(\req_msg[6] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U9 ( .Z(\dpath/b_mux_out[7] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[7] ), .A2(\req_msg[7] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U10 ( .Z(\dpath/b_mux_out[8] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[8] ), .A2(\req_msg[8] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U11 ( .Z(\dpath/b_mux_out[9] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[9] ), .A2(\req_msg[9] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U12 ( .Z(\dpath/b_mux_out[10] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[10] ), .A2(\req_msg[10] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U13 ( .Z(\dpath/b_mux_out[11] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[11] ), .A2(\req_msg[11] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U14 ( .Z(\dpath/b_mux_out[12] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[12] ), .A2(\req_msg[12] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U15 ( .Z(\dpath/b_mux_out[13] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[13] ), .A2(\req_msg[13] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U16 ( .Z(\dpath/b_mux_out[14] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[14] ), .A2(\req_msg[14] ), .A1(ctrl_b_mux_sel_0_ ) );
AO22D1BWP40P140 \dpath/b_mux/U17 ( .Z(\dpath/b_mux_out[15] ), .B2(\dpath/b_mux/n1 ), .B1(\dpath/a_reg_out[15] ), .A2(\req_msg[15] ), .A1(ctrl_b_mux_sel_0_ ) );
INVD3BWP40P140 \dpath/sub/U1 ( .ZN(\resp_msg[1] ), .I(\dpath/sub/n1 ) );
INVD3BWP40P140 \dpath/sub/U2 ( .ZN(\resp_msg[11] ), .I(\dpath/sub/n11 ) );
INVD3BWP40P140 \dpath/sub/U3 ( .ZN(\resp_msg[12] ), .I(\dpath/sub/n9 ) );
INVD3BWP40P140 \dpath/sub/U4 ( .ZN(\resp_msg[13] ), .I(\dpath/sub/n7 ) );
INVD3BWP40P140 \dpath/sub/U5 ( .ZN(\resp_msg[14] ), .I(\dpath/sub/n5 ) );
INVD3BWP40P140 \dpath/sub/U6 ( .ZN(\resp_msg[6] ), .I(\dpath/sub/n3 ) );
INVD1BWP40P140 \dpath/sub/U7 ( .ZN(\dpath/sub/n44 ), .I(\dpath/b_reg_out[0] ) );
INVD1BWP40P140 \dpath/sub/U8 ( .ZN(\dpath/sub/n5 ), .I(\dpath/sub/n45 ) );
INVD1BWP40P140 \dpath/sub/U9 ( .ZN(\dpath/sub/n7 ), .I(\dpath/sub/n46 ) );
INVD1BWP40P140 \dpath/sub/U10 ( .ZN(\dpath/sub/n9 ), .I(\dpath/sub/n47 ) );
INVD1BWP40P140 \dpath/sub/U11 ( .ZN(\dpath/sub/n11 ), .I(\dpath/sub/n48 ) );
FA1D4BWP40P140 \dpath/sub/U12 ( .S(\resp_msg[10] ), .CO(\dpath/sub/n27 ), .CI(\dpath/sub/n19 ), .B(\dpath/sub/n20 ), .A(\dpath/a_reg_out[10] ) );
FA1D4BWP40P140 \dpath/sub/U13 ( .S(\resp_msg[9] ), .CO(\dpath/sub/n19 ), .CI(\dpath/sub/n29 ), .B(\dpath/a_reg_out[9] ), .A(\dpath/sub/n30 ) );
FA1D4BWP40P140 \dpath/sub/U14 ( .S(\resp_msg[8] ), .CO(\dpath/sub/n29 ), .CI(\dpath/sub/n21 ), .B(\dpath/a_reg_out[8] ), .A(\dpath/sub/n22 ) );
FA1D4BWP40P140 \dpath/sub/U15 ( .S(\resp_msg[7] ), .CO(\dpath/sub/n21 ), .CI(\dpath/sub/n31 ), .B(\dpath/a_reg_out[7] ), .A(\dpath/sub/n32 ) );
FA1D4BWP40P140 \dpath/sub/U16 ( .S(\resp_msg[5] ), .CO(\dpath/sub/n23 ), .CI(\dpath/sub/n33 ), .B(\dpath/sub/n34 ), .A(\dpath/a_reg_out[5] ) );
FA1D4BWP40P140 \dpath/sub/U17 ( .S(\resp_msg[4] ), .CO(\dpath/sub/n33 ), .CI(\dpath/sub/n25 ), .B(\dpath/a_reg_out[4] ), .A(\dpath/sub/n26 ) );
FA1D4BWP40P140 \dpath/sub/U18 ( .S(\resp_msg[3] ), .CO(\dpath/sub/n25 ), .CI(\dpath/sub/n35 ), .B(\dpath/a_reg_out[3] ), .A(\dpath/sub/n36 ) );
FA1D4BWP40P140 \dpath/sub/U19 ( .S(\resp_msg[2] ), .CO(\dpath/sub/n35 ), .CI(\dpath/sub/n15 ), .B(\dpath/a_reg_out[2] ), .A(\dpath/sub/n16 ) );
OR2D1BWP40P140 \dpath/sub/U20 ( .Z(\dpath/sub/n13 ), .A2(\dpath/a_reg_out[0] ), .A1(\dpath/sub/n44 ) );
INVD1BWP40P140 \dpath/sub/U21 ( .ZN(\dpath/sub/n20 ), .I(\dpath/b_reg_out[10] ) );
INVD1BWP40P140 \dpath/sub/U22 ( .ZN(\dpath/sub/n28 ), .I(\dpath/b_reg_out[11] ) );
INVD1BWP40P140 \dpath/sub/U23 ( .ZN(\dpath/sub/n32 ), .I(\dpath/b_reg_out[7] ) );
INVD1BWP40P140 \dpath/sub/U24 ( .ZN(\dpath/sub/n30 ), .I(\dpath/b_reg_out[9] ) );
INVD1BWP40P140 \dpath/sub/U25 ( .ZN(\dpath/sub/n24 ), .I(\dpath/b_reg_out[6] ) );
INVD1BWP40P140 \dpath/sub/U26 ( .ZN(\dpath/sub/n36 ), .I(\dpath/b_reg_out[3] ) );
INVD1BWP40P140 \dpath/sub/U27 ( .ZN(\dpath/sub/n26 ), .I(\dpath/b_reg_out[4] ) );
INVD1BWP40P140 \dpath/sub/U28 ( .ZN(\dpath/sub/n34 ), .I(\dpath/b_reg_out[5] ) );
INVD1BWP40P140 \dpath/sub/U29 ( .ZN(\dpath/sub/n14 ), .I(\dpath/b_reg_out[1] ) );
INVD1BWP40P140 \dpath/sub/U30 ( .ZN(\dpath/sub/n16 ), .I(\dpath/b_reg_out[2] ) );
FA1D1BWP40P140 \dpath/sub/U31 ( .S(\dpath/sub/n49 ), .CO(\dpath/sub/n31 ), .CI(\dpath/sub/n23 ), .B(\dpath/a_reg_out[6] ), .A(\dpath/sub/n24 ) );
FA1D1BWP40P140 \dpath/sub/U32 ( .S(\dpath/sub/n48 ), .CO(\dpath/sub/n17 ), .CI(\dpath/sub/n27 ), .B(\dpath/a_reg_out[11] ), .A(\dpath/sub/n28 ) );
FA1D1BWP40P140 \dpath/sub/U33 ( .S(\dpath/sub/n45 ), .CO(\dpath/sub/n42 ), .CI(\dpath/sub/n40 ), .B(\dpath/a_reg_out[14] ), .A(\dpath/sub/n41 ) );
INVD1BWP40P140 \dpath/sub/U34 ( .ZN(\dpath/sub/n41 ), .I(\dpath/b_reg_out[14] ) );
FA1D1BWP40P140 \dpath/sub/U35 ( .S(\dpath/sub/n50 ), .CO(\dpath/sub/n15 ), .CI(\dpath/sub/n13 ), .B(\dpath/a_reg_out[1] ), .A(\dpath/sub/n14 ) );
FA1D1BWP40P140 \dpath/sub/U36 ( .S(\dpath/sub/n47 ), .CO(\dpath/sub/n37 ), .CI(\dpath/sub/n17 ), .B(\dpath/a_reg_out[12] ), .A(\dpath/sub/n18 ) );
INVD1BWP40P140 \dpath/sub/U37 ( .ZN(\dpath/sub/n18 ), .I(\dpath/b_reg_out[12] ) );
FA1D1BWP40P140 \dpath/sub/U38 ( .S(\dpath/sub/n46 ), .CO(\dpath/sub/n40 ), .CI(\dpath/sub/n37 ), .B(\dpath/a_reg_out[13] ), .A(\dpath/sub/n38 ) );
INVD1BWP40P140 \dpath/sub/U39 ( .ZN(\dpath/sub/n38 ), .I(\dpath/b_reg_out[13] ) );
XNR2UD1BWP40P140 \dpath/sub/U40 ( .ZN(\dpath/n15 ), .A2(\dpath/sub/n44 ), .A1(\dpath/a_reg_out[0] ) );
INVD1BWP40P140 \dpath/sub/U41 ( .ZN(\dpath/sub/n1 ), .I(\dpath/sub/n50 ) );
INVD1BWP40P140 \dpath/sub/U42 ( .ZN(\dpath/sub/n3 ), .I(\dpath/sub/n49 ) );
XOR2UD1BWP40P140 \dpath/sub/U43 ( .Z(\dpath/sub/n43 ), .A2(\dpath/a_reg_out[15] ), .A1(\dpath/sub/n39 ) );
INVD1BWP40P140 \dpath/sub/U44 ( .ZN(\dpath/sub/n22 ), .I(\dpath/b_reg_out[8] ) );
INVD1BWP40P140 \dpath/sub/U45 ( .ZN(\dpath/sub/n39 ), .I(\dpath/b_reg_out[15] ) );
XOR2D4BWP40P140 \dpath/sub/U46 ( .Z(\resp_msg[15] ), .A2(\dpath/sub/n42 ), .A1(\dpath/sub/n43 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_15_ ( .Q(\dpath/b_reg_out[15] ), .D(\dpath/b_reg/n17 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_14_ ( .Q(\dpath/b_reg_out[14] ), .D(\dpath/b_reg/n16 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_13_ ( .Q(\dpath/b_reg_out[13] ), .D(\dpath/b_reg/n15 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_12_ ( .Q(\dpath/b_reg_out[12] ), .D(\dpath/b_reg/n14 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_11_ ( .Q(\dpath/b_reg_out[11] ), .D(\dpath/b_reg/n13 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_10_ ( .Q(\dpath/b_reg_out[10] ), .D(\dpath/b_reg/n12 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_9_ ( .Q(\dpath/b_reg_out[9] ), .D(\dpath/b_reg/n11 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_8_ ( .Q(\dpath/b_reg_out[8] ), .D(\dpath/b_reg/n10 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_7_ ( .Q(\dpath/b_reg_out[7] ), .D(\dpath/b_reg/n9 ), .CP(clk_1 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_6_ ( .Q(\dpath/b_reg_out[6] ), .D(\dpath/b_reg/n8 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_5_ ( .Q(\dpath/b_reg_out[5] ), .D(\dpath/b_reg/n7 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_4_ ( .Q(\dpath/b_reg_out[4] ), .D(\dpath/b_reg/n6 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_3_ ( .Q(\dpath/b_reg_out[3] ), .D(\dpath/b_reg/n5 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_2_ ( .Q(\dpath/b_reg_out[2] ), .D(\dpath/b_reg/n4 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_0_ ( .Q(\dpath/b_reg_out[0] ), .D(\dpath/b_reg/n2 ), .CP(clk_0 ) );
DFQD1BWP40P140 \dpath/b_reg/out_reg_1_ ( .Q(\dpath/b_reg_out[1] ), .D(\dpath/b_reg/n3 ), .CP(clk_0 ) );
INVD1BWP40P140 \dpath/b_reg/U2 ( .ZN(\dpath/b_reg/n1 ), .I(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U3 ( .Z(\dpath/b_reg/n17 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[15] ), .A2(\dpath/b_mux_out[15] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U4 ( .Z(\dpath/b_reg/n16 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[14] ), .A2(\dpath/b_mux_out[14] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U5 ( .Z(\dpath/b_reg/n15 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[13] ), .A2(\dpath/b_mux_out[13] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U6 ( .Z(\dpath/b_reg/n14 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[12] ), .A2(\dpath/b_mux_out[12] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U7 ( .Z(\dpath/b_reg/n13 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[11] ), .A2(\dpath/b_mux_out[11] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U8 ( .Z(\dpath/b_reg/n12 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[10] ), .A2(\dpath/b_mux_out[10] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U9 ( .Z(\dpath/b_reg/n11 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[9] ), .A2(\dpath/b_mux_out[9] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U10 ( .Z(\dpath/b_reg/n10 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[8] ), .A2(\dpath/b_mux_out[8] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U11 ( .Z(\dpath/b_reg/n9 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[7] ), .A2(\dpath/b_mux_out[7] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U12 ( .Z(\dpath/b_reg/n8 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[6] ), .A2(\dpath/b_mux_out[6] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U13 ( .Z(\dpath/b_reg/n7 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[5] ), .A2(\dpath/b_mux_out[5] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U14 ( .Z(\dpath/b_reg/n6 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[4] ), .A2(\dpath/b_mux_out[4] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U15 ( .Z(\dpath/b_reg/n5 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[3] ), .A2(\dpath/b_mux_out[3] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U16 ( .Z(\dpath/b_reg/n4 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[2] ), .A2(\dpath/b_mux_out[2] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U17 ( .Z(\dpath/b_reg/n3 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[1] ), .A2(\dpath/b_mux_out[1] ), .A1(ctrl_b_reg_en_0_ ) );
AO22D1BWP40P140 \dpath/b_reg/U18 ( .Z(\dpath/b_reg/n2 ), .B2(\dpath/b_reg/n1 ), .B1(\dpath/b_reg_out[0] ), .A2(\dpath/b_mux_out[0] ), .A1(ctrl_b_reg_en_0_ ) );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_1 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_2 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_3 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_4 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_5 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_6 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_7 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_8 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_9 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_10 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_11 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_12 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_13 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_14 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_15 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_16 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_17 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_18 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_19 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_20 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_21 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_22 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_23 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_24 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_25 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_26 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_27 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_28 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_29 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_30 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_31 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_32 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_33 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_34 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_35 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_36 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_37 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_38 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_39 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_40 (  );
BOUNDARY_LEFTBWP40P140 BNDRY_CAP_41 (  );
BOUNDARY_RIGHTBWP40P140 BNDRY_CAP_42 (  );
TAPCELLBWP40P140 WELLTAP_1 (  );
TAPCELLBWP40P140 WELLTAP_2 (  );
TAPCELLBWP40P140 WELLTAP_3 (  );
TAPCELLBWP40P140 WELLTAP_4 (  );
TAPCELLBWP40P140 WELLTAP_5 (  );
TAPCELLBWP40P140 WELLTAP_6 (  );
TAPCELLBWP40P140 WELLTAP_7 (  );
TAPCELLBWP40P140 WELLTAP_8 (  );
TAPCELLBWP40P140 WELLTAP_9 (  );
TAPCELLBWP40P140 WELLTAP_10 (  );
TAPCELLBWP40P140 WELLTAP_11 (  );
TAPCELLBWP40P140 WELLTAP_12 (  );
TAPCELLBWP40P140 WELLTAP_13 (  );
TAPCELLBWP40P140 WELLTAP_14 (  );
TAPCELLBWP40P140 WELLTAP_15 (  );
TAPCELLBWP40P140 WELLTAP_16 (  );
TAPCELLBWP40P140 WELLTAP_17 (  );
TAPCELLBWP40P140 WELLTAP_18 (  );
TAPCELLBWP40P140 WELLTAP_19 (  );
TAPCELLBWP40P140 WELLTAP_20 (  );
TAPCELLBWP40P140 WELLTAP_21 (  );
TAPCELLBWP40P140 WELLTAP_22 (  );
TAPCELLBWP40P140 WELLTAP_23 (  );
DCAP4BWP40P140 BNDRY_CAP_TAP_1 (  );
DCAP4BWP40P140 BNDRY_CAP_TAP_2 (  );
DCAP64BWP40P140HVT BNDRY_CAP_43 (  );
DCAP32BWP40P140HVT BNDRY_CAP_44 (  );
DCAP16BWP40P140HVT BNDRY_CAP_45 (  );
DCAP4BWP40P140HVT BNDRY_CAP_46 (  );
FILL2BWP40P140HVT BNDRY_CAP_47 (  );
DCAP64BWP40P140HVT BNDRY_CAP_48 (  );
DCAP32BWP40P140HVT BNDRY_CAP_49 (  );
DCAP16BWP40P140HVT BNDRY_CAP_50 (  );
DCAP4BWP40P140HVT BNDRY_CAP_51 (  );
FILL2BWP40P140HVT BNDRY_CAP_52 (  );
BUFFD3BWP30P140LVT clk_0_buf ( .Z(clk_0 ), .I(clk ) );
BUFFD4BWP30P140LVT clk_1_buf ( .Z(clk_1 ), .I(clk ) );

endmodule
